leon.fuchs@tallinn.emse.fr.209947:1702021731