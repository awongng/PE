//Name of file
//Description of module behavior

`timescale 1ps/1ns

module module_name (
    input logic [31:0] input_example_i;
    input logic input_example_2_i
    output logic [31:0] output_example_o;
);
    logic



endmodule:module_name